import(<kernel.cdl>);

/* mrubyの本体 */
import(<tMruby.cdl>);

import("sMrubyUDP.cdl");
import("sMrubyTCP.cdl");

/*
 * シグニチャプラグイン MrubyBridgePlugin の呼び出し。
 */
generate( MrubyBridgePlugin, sKernel, "" );
generate( MrubyBridgePlugin, sMrubyUDP, "" );
generate( MrubyBridgePlugin, sMrubyTCP, "" );

/*
 *  サンプルプログラムの定義
 */
cell nMruby::tsKernel BridgeKernel {
	cTECS = Kernel.eKernel;
};

cell nMruby::tsMrubyUDP BridgeUDP {
	cTECS = MrubyUDP.eMrubyUDP;
};

cell nMruby::tsMrubyTCP BridgeTCP {
	cTECS = MrubyTCP.eMrubyTCP;
};

cell tMrubyUDP MrubyUDP {
	cAPI = UDPCEP_000.eAPI;
};

cell tMrubyTCP MrubyTCP {
	cAPI = TCPCEP_000.eAPI;
	cREP4_000 = REP4_000.eREP4;
    cRepSelector = RepSelector.eRepSelector;
};