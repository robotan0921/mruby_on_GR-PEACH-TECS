import(<bridge.cdl>);

cell nMruby::tMruby Mruby {
	mrubyFile =
		"$(MRUBY_LIB_DIR)/RTOS.rb "
		"$(MRUBY_LIB_DIR)/LED.rb "
		"$(MRUBY_APP_DIR)/led_sample.rb";

	cInit = VM_TECSInitializer.eInitialize;
    cSerialPort = SerialPort1.eSerialPort;
};

cell tTask MrubyTask1 {
	cTaskBody = Mruby.eMrubyBody;
	attribute = C_EXP("TA_ACT");
	priority  = 10;
    stackSize = 4096;
};
