import(<kernel.cdl>);

/* mrubyの本体 */
import(<tMruby.cdl>);

import(<tLED.cdl>);

/*
 * シグニチャプラグイン MrubyBridgePlugin の呼び出し。
 */
generate( MrubyBridgePlugin, sKernel, "" );
generate( MrubyBridgePlugin, sLED, "" );

/*
 *  サンプルプログラムの定義
 */
cell nMruby::tsKernel BridgeKernel {
	cTECS = Kernel.eKernel;
};
cell nMruby::tsLED BridgeLED {
	cTECS = LED.eLED;
};


cell tLED LED {};
