signature sMrubyUDP {
    ER_UINT send([in,size_is(len)]const char_t *data, [in]int32_t len, [in]uint32_t dstaddr,
                 [in]uint16_t dstport, [in]TMO tmout);
    ER_UINT receive([out,size_is(len)]char_t *data, [in]int32_t len, [in]TMO tmout);
    ER cancelSend([in]ER error);
    ER cancelReceive([in]ER error);

    uint32_t make_ipv4_addr([in]uint32_t a, [in]uint32_t b, [in]uint32_t c, [in]uint32_t d);
};

celltype tMrubyUDP {
    call sUDPCEPAPI4 cAPI;
	entry sMrubyUDP eMrubyUDP;
};