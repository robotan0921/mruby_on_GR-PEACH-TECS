
[singleton, active]
celltype tIfMbedAdapter {
	call	sNicDriver cNicDriver;
};