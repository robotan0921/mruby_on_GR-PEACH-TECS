/*
 *		C言語で記述されたアプリケーションから，TECSベースの実行時間分布
 *		集計サービスを呼び出すためのアダプタ用セルタイプの定義
 * 
 *  $Id: tHistogramAdapter.cdl 509 2016-01-12 06:06:14Z ertl-hiro $
 */
[singleton, active]
celltype tHistogramAdapter {
	call	sHistogram		cHistogram[];
};
