signature sMrubyTCP {
    ER      accept([in]uint16_t descid, [out]uint32_t *ipaddr, [out]uint16_t *portno, [in]TMO tmout);
    ER      connect([in]T_IN4_ADDR myaddr, [in]uint16_t myport, [in]T_IN4_ADDR dstaddr, [in]uint16_t dstport, [in]TMO tmout);
    ER_UINT send([in,size_is(len)]const char_t *data, [in]int32_t len, [in]TMO tmout);
    ER_UINT receive([out,size_is(len)]char_t *data, [in]int32_t len, [in]TMO tmout);
    ER      cancel([in]FN fncd);
    ER      close([in]TMO tmout);
    ER      shutdown(void);

    uint32_t make_ipv4_addr([in]uint32_t a, [in]uint32_t b, [in]uint32_t c, [in]uint32_t d);
};

celltype tMrubyTCP {
    call sTCPCEPAPI4 cAPI;
	call sREP4 cREP4_000;
    call sRepSelector cRepSelector;

	entry sMrubyTCP eMrubyTCP;
};