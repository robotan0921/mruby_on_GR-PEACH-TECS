import(<kernel.cdl>);

/* mrubyの本体 */
import(<tMruby.cdl>);

import(<tLED.cdl>);
import(<tButton.cdl>);


/*
 * シグニチャプラグイン MrubyBridgePlugin の呼び出し。
 */
generate( MrubyBridgePlugin, sKernel, "" );
generate( MrubyBridgePlugin, sLED, "" );
generate( MrubyBridgePlugin, sButton, "" );

/*
 *  サンプルプログラムの定義
 */
cell nMruby::tsKernel BridgeKernel {
	cTECS = Kernel.eKernel;
};
cell nMruby::tsLED BridgeLED {
	cTECS = LED.eLED;
};
cell nMruby::tsButton BridgeButton {
	cTECS = Button.eButton;
};


cell tLED LED {};
cell tButton Button {};
